
(* Exercise 8.3
Define the reflexive and transitive closure of a binary relation
(using an inductive definition). The Rstar module of the Coq
standard library provides an impredicative definition of this
closure (constant Rstar). Prove that the two definitions are equal.
*)